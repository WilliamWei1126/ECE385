`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/16/2026 10:51:29 PM
// Design Name: 
// Module Name: 9BitAdder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NineBitAdder(
    input logic[8:0] In1,
    input logic[8:0] In2,
    
    output logic[8:0] Result
    );
endmodule
