module ece385_gnd(
        output logic GND
    );
    
    assign GND = 1'b0; // What did you expect?
    
endmodule
